module OBUF (
    output logic O,
    input  logic I
);
    assign O = I;
endmodule // OBUF
