module IBUF (
    output logic O,
    input  logic I
);
    assign O = I;
endmodule // IBUF
